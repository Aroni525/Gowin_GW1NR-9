module Global;

integer CrystalClockMhz = 27;

endmodule